library verilog;
use verilog.vl_types.all;
entity dividable11_vlg_vec_tst is
end dividable11_vlg_vec_tst;
