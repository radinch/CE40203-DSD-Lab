library verilog;
use verilog.vl_types.all;
entity Compare_4_vlg_vec_tst is
end Compare_4_vlg_vec_tst;
