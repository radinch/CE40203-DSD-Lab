library verilog;
use verilog.vl_types.all;
entity divideable3_vlg_vec_tst is
end divideable3_vlg_vec_tst;
