library verilog;
use verilog.vl_types.all;
entity dividable11_vlg_check_tst is
    port(
        ans             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end dividable11_vlg_check_tst;
