library verilog;
use verilog.vl_types.all;
entity waitingRoom_vlg_vec_tst is
end waitingRoom_vlg_vec_tst;
