module tb;
    reg [3:0] A;
    reg [3:0] B;
    wire lt, gt, eq;

    // Instantiate the 4-bit comparator
    FourBitComparator uut (
        .A(A),
        .B(B),
        .lt(lt),
        .gt(gt),
        .eq(eq)
    );

    initial begin
        // Monitor the changes in A, B, lt, gt, eq
        $monitor("A = %b, B = %b, lt = %b, gt = %b, eq = %b", A, B, lt, gt, eq);
        
        // Test all possible combinations
        A = 4'b0000; B = 4'b0000; #10;
        A = 4'b0001; B = 4'b0000; #10;
        A = 4'b0001; B = 4'b0001; #10;
        A = 4'b0010; B = 4'b0001; #10;
        A = 4'b0011; B = 4'b0001; #10;
        A = 4'b0100; B = 4'b0001; #10;
        A = 4'b0101; B = 4'b0001; #10;
        A = 4'b0110; B = 4'b0001; #10;
        A = 4'b0111; B = 4'b0001; #10;
        A = 4'b1000; B = 4'b0001; #10;
        A = 4'b1001; B = 4'b0001; #10;
        A = 4'b1010; B = 4'b0001; #10;
        A = 4'b1011; B = 4'b0001; #10;
        A = 4'b1100; B = 4'b0001; #10;
        A = 4'b1101; B = 4'b0001; #10;
        A = 4'b1110; B = 4'b0001; #10;
        A = 4'b1111; B = 4'b0001; #10;

        // Test all combinations where A is less than B
        A = 4'b0000; B = 4'b0001; #10;
        A = 4'b0000; B = 4'b0010; #10;
        A = 4'b0000; B = 4'b0011; #10;
        A = 4'b0000; B = 4'b0100; #10;
        A = 4'b0000; B = 4'b0101; #10;
        A = 4'b0000; B = 4'b0110; #10;
        A = 4'b0000; B = 4'b0111; #10;
        A = 4'b0000; B = 4'b1000; #10;
        A = 4'b0000; B = 4'b1001; #10;
        A = 4'b0000; B = 4'b1010; #10;
        A = 4'b0000; B = 4'b1011; #10;
        A = 4'b0000; B = 4'b1100; #10;
        A = 4'b0000; B = 4'b1101; #10;
        A = 4'b0000; B = 4'b1110; #10;
        A = 4'b0000; B = 4'b1111; #10;

        // Test all combinations where A is greater than B
        A = 4'b0001; B = 4'b0000; #10;
        A = 4'b0010; B = 4'b0000; #10;
        A = 4'b0011; B = 4'b0000; #10;
        A = 4'b0100; B = 4'b0000; #10;
        A = 4'b0101; B = 4'b0000; #10;
        A = 4'b0110; B = 4'b0000; #10;
        A = 4'b0111; B = 4'b0000; #10;
        A = 4'b1000; B = 4'b0000; #10;
        A = 4'b1001; B = 4'b0000; #10;
        A = 4'b1010; B = 4'b0000; #10;
        A = 4'b1011; B = 4'b0000; #10;
        A = 4'b1100; B = 4'b0000; #10;
        A = 4'b1101; B = 4'b0000; #10;
        A = 4'b1110; B = 4'b0000; #10;
        A = 4'b1111; B = 4'b0000; #10;

        // Test all combinations where A is equal to B
        A = 4'b0000; B = 4'b0000; #10;
        A = 4'b0001; B = 4'b0001; #10;
        A = 4'b0010; B = 4'b0010; #10;
        A = 4'b0011; B = 4'b0011; #10;
        A = 4'b0100; B = 4'b0100; #10;
        A = 4'b0101; B = 4'b0101; #10;
        A = 4'b0110; B = 4'b0110; #10;
        A = 4'b0111; B = 4'b0111; #10;
        A = 4'b1000; B = 4'b1000; #10;
        A = 4'b1001; B = 4'b1001; #10;
        A = 4'b1010; B = 4'b1010; #10;
        A = 4'b1011; B = 4'b1011; #10;
        A = 4'b1100; B = 4'b1100; #10;
        A = 4'b1101; B = 4'b1101; #10;
        A = 4'b1110; B = 4'b1110; #10;
        A = 4'b1111; B = 4'b1111; #10;
        
        $stop;
    end
endmodule
