library verilog;
use verilog.vl_types.all;
entity Compare_2_vlg_vec_tst is
end Compare_2_vlg_vec_tst;
